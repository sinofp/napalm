module fetch (/*AUTOARG*/ ) ;
   
endmodule // fetch
