module decode (/*AUTOARG*/ ) ;
   
endmodule // decode
