`timescale 1ns / 1ps

module reg_heap (
    input[4:0] ra1,
    input[4:0] ra2,
    input[4:0] wa,
    input we,
    input[31:0] wd,
    output[31:0] rd1,
    output[31:0] rd2
);
    
endmodule