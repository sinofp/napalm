module writeback (/*AUTOARG*/ ) ;
   
endmodule // writeback
