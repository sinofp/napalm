`timescale 1ns / 1ps

module data_mem (
         input[31:0] addr, // TODO
         input[31:0] wd,
         input we,
         output[31:0] rd
       );

endmodule
