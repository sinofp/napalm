module memory (/*AUTOARG*/ ) ;
   
endmodule // memory
