module alu (
           input[5:0] op_code,
           input[31:0] num1,
           input[31:0] num2,
           output[31:0] res
       );

endmodule
